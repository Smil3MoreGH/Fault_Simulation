// IWLS benchmark module "C17.iscas" printed on Wed Mar  6 23:40:18 2002

module \C17.iscas ( 
    \1GAT(0) , \2GAT(1) ,\22GAT(10) );
    
  input  \1GAT(0), \2GAT(1) ;
  output \22GAT(10) ;
  
  assign \22GAT(10)  = \1GAT(0)  | \2GAT(1) ;

endmodule
